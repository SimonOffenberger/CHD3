-------------------------------------------------------------------------------
-- Title : PosEdgeTrigDFF
-- Project : Chip Design 3
-------------------------------------------------------------------------------
-- File : PosEdgeTrigDFF-AsyncSeq-a.vhd
-- Author : 
-- Created : 2006-11-05
-- Last update: 2012-11-21
-------------------------------------------------------------------------------
-- Copyright (c) Hagenberg/Austria 2006-2012
-------------------------------------------------------------------------------
-- Subversion entries:
-- $Id: $
-------------------------------------------------------------------------------
-- Description:
-- Implementation of a positive edge triggered D-FF based on trational 
-- NAND gates.
-------------------------------------------------------------------------------

architecture AsyncSeq of PosEdgeTrigDFF is

begin  -- AsyncSeq

  ---------------------------------------------------------------------------------------
  -- Add your code here
  ---------------------------------------------------------------------------------------

end AsyncSeq;
