library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.global.all;

entity tbMultiplier is
end tbMultiplier;


architecture Bhv of tbMultiplier is

  -- ------------------------------------------------------
  -- add your code here (signal, constant, ... declaration)
  -- ------------------------------------------------------

begin
  
  -- ------------------
  -- add your code here
  -- ------------------

  -- Test loop for multiplicant and multiplier to verify completeness
  TestSequence : process is
  begin
  
  -- ------------------
  -- add your code here
  -- ------------------

  end process TestSequence;
  
end Bhv;

