-------------------------------------------------------------------------------
-- Title : Sync Stage
-- Project : Chip Design
-------------------------------------------------------------------------------
-- Author : simon Offenberger
-- Created : 2025-12-1
-------------------------------------------------------------------------------
-- Copyright (c) Hagenberg/Austria 2015
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Entity 
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity EdgeDetection is
  port (
    iClk : in std_ulogic;
    inResetAsync : in std_ulogic;
    iEnable : in std_ulogic;
    iSync : in std_ulogic;
    oEdge : out std_ulogic);
end EdgeDetection;