-------------------------------------------------------------------------------
-- Title : Running Light
-- Project : Chip Design
-------------------------------------------------------------------------------
-- Author : simon Offenberger
-- Created : 2025-11-11
-------------------------------------------------------------------------------
-- Copyright (c) Hagenberg/Austria 2015
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Entity 
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity RunningLight is
 port (
  iClk         : in std_ulogic;
  inResetAsync : in std_ulogic;
  iEnable      : in std_ulogic;
  oState       : out std_ulogic_vector(2 downto 0));
 end RunningLight;
