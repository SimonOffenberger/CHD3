---------------------------------------------------------------------------
-- Title      : Testbench for HelloDE1
-- Project    : HelloDE1
-- Company    : FH OOe Hagenberg/A, Copyright (c) 2015
-------------------------------------------------------------------------------
-- Author	  : Thomas Mueller-W,
-- Date		  : 30.4.2015
-- Authors are
-- 		tm	  : Thomas Mueller-W., Hagenberg
-- Revisions  : V1, 30.4.15, tm
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity tbHello is
end tbHello;
